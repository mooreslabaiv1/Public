


class weighted_round_robin_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_test extends weighted_round_robin_base_test;

  `uvm_component_utils(weighted_round_robin_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_test)

  function new(string name="weighted_round_robin_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_test", uvm_component parent=null);
    super.new(name, parent);
  endfunction

  virtual task run_phase(uvm_phase phase);
    // Declarations at the beginning of the task as per coding guidelines
    rr_request_seq_pkg::rr_request_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_sequence m_rr_request_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq;
    rr_grant_monitor_seq_pkg::rr_grant_monitor_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_sequence m_rr_grant_monitor_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq;
    prio_update_seq_pkg::prio_update_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_sequence m_prio_update_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq;

    super.run_phase(phase);
    phase.raise_objection(this);

    // Create sequences prior to fork as required
    m_rr_request_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq =
      rr_request_seq_pkg::rr_request_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_sequence::type_id::create("m_rr_request_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq");
    m_rr_grant_monitor_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq =
      rr_grant_monitor_seq_pkg::rr_grant_monitor_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_sequence::type_id::create("m_rr_grant_monitor_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq");
    m_prio_update_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq =
      prio_update_seq_pkg::prio_update_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_sequence::type_id::create("m_prio_update_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq");

    fork
      m_rr_request_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq.start(m_env.m_rr_request_agent.m_seqr);
      m_rr_grant_monitor_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq.start(m_env.m_rr_grant_monitor_agent.m_seqr);
      m_prio_update_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_seq.start(m_env.m_prio_update_agent.m_seqr);
    join_any

    phase.drop_objection(this);
  endtask

endclass : weighted_round_robin_arbiter_maximal_concurrent_requests_and_dynamic_priority_update_stress_test_test