package wrr_arbitration_seq_pkg;

  //******************************************************************************
  // Imports
  //******************************************************************************
  import uvm_pkg::*;
  import wrr_arbitration_agent_pkg::*;
  `include "uvm_macros.svh"

  //******************************************************************************
  // Includes
  //******************************************************************************
  `include "wrr_arbitration_base_seq.sv"

endpackage : wrr_arbitration_seq_pkg