


    `ifndef FSM_SEEK_DETECT_ENV_INC_SV
    `define FSM_SEEK_DETECT_ENV_INC_SV
    `include "tb_src.incl"    
    `include "fsm_seek_detect_env_cfg.sv"
    // Include the reference model here
    `include "fsm_seek_detect_ref_model.sv"

    `include "fsm_seek_detect_sbd.sv"
    
    `include "fsm_seek_detect_fsm_seek_detect_monitor_env_cov.sv"
    `include "fsm_seek_detect_fsm_seek_detect_monitor_connect_cov.sv"


    // <Optional> ToDo: Add additional required `include directives
    
    `endif // FSM_SEEK_DETECT_ENV_INC_SV
    