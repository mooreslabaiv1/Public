package requestor_seq_pkg;

    //******************************************************************************
    // Imports
    //******************************************************************************
    import uvm_pkg::*;
    import requestor_agent_pkg::*;

    //******************************************************************************
    // Includes
    //******************************************************************************
    `include "requestor_base_seq.sv"
    `include "requestor_basic_functionality_seq.sv"

endpackage : requestor_seq_pkg
