package prio_update_agent_pkg;

  //******************************************************************************
  // Imports
  //******************************************************************************
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  //******************************************************************************
  // Includes
  //******************************************************************************
  `include "prio_update_trans_item.sv"
  `include "prio_update_monitor.sv"
  `include "prio_update_driver.sv"
  `include "prio_update_seqr.sv"
  `include "prio_update_agent_cov.sv"
  `include "prio_update_agent_cfg.sv"
  `include "prio_update_agent.sv"

endpackage : prio_update_agent_pkg