
package rr_grant_monitor_agent_pkg;

  //******************************************************************************
  // Imports
  //******************************************************************************
  import uvm_pkg::*;

  //******************************************************************************
  // Includes
  //******************************************************************************
  `include "rr_grant_monitor_trans_item.sv"
  `include "rr_grant_monitor_monitor.sv"
  `include "rr_grant_monitor_driver.sv"
  `include "rr_grant_monitor_seqr.sv"
  `include "rr_grant_monitor_agent_cov.sv"
  `include "rr_grant_monitor_agent_cfg.sv"
  `include "rr_grant_monitor_agent.sv"

endpackage : rr_grant_monitor_agent_pkg