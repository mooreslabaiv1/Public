package prio_update_seq_pkg;

    //******************************************************************************
    // Imports
    //******************************************************************************
    import uvm_pkg::*;
    import prio_update_agent_pkg::*;

    //******************************************************************************
    // Includes
    //******************************************************************************
    `include "prio_update_base_seq.sv"
    `include "prio_update_basic_functionality_seq.sv"

endpackage : prio_update_seq_pkg
