package wrr_prio_update_agent_pkg;

  //******************************************************************************
  // Imports
  //******************************************************************************
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  //******************************************************************************
  // Includes
  //******************************************************************************
  `include "wrr_prio_update_trans_item.sv"
  `include "wrr_prio_update_monitor.sv"
  `include "wrr_prio_update_driver.sv"
  `include "wrr_prio_update_seqr.sv"
  `include "wrr_prio_update_agent_cov.sv"
  `include "wrr_prio_update_agent_cfg.sv"
  `include "wrr_prio_update_agent.sv"

endpackage : wrr_prio_update_agent_pkg