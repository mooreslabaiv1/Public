package serial_agent_pkg;

  //******************************************************************************
  // Imports
  //******************************************************************************
  import uvm_pkg::*;

  //******************************************************************************
  // Includes
  //******************************************************************************
  `include "serial_trans_item.sv"
  `include "serial_monitor.sv"
  `include "serial_driver.sv"
  `include "serial_seqr.sv"
  `include "serial_agent_cov.sv"
  `include "serial_agent_cfg.sv"
  `include "serial_agent.sv"

endpackage : serial_agent_pkg