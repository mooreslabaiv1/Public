package wrr_prio_update_seq_pkg;

  //******************************************************************************
  // Imports
  //******************************************************************************
  import uvm_pkg::*;
  import wrr_prio_update_agent_pkg::*;
  `include "uvm_macros.svh"

  //******************************************************************************
  // Includes
  //******************************************************************************
  `include "wrr_prio_update_base_seq.sv"

endpackage : wrr_prio_update_seq_pkg