package rr_request_agent_pkg;

  //******************************************************************************
  // Imports
  //******************************************************************************
  import uvm_pkg::*;

  //******************************************************************************
  // Includes
  //******************************************************************************
  `include "rr_request_trans_item.sv"
  `include "rr_request_monitor.sv"
  `include "rr_request_driver.sv"
  `include "rr_request_seqr.sv"
  `include "rr_request_agent_cov.sv"
  `include "rr_request_agent_cfg.sv"
  `include "rr_request_agent.sv"

endpackage : rr_request_agent_pkg