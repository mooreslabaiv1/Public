package clk_rst_seq_pkg;

  //******************************************************************************
  // Imports
  //******************************************************************************
  import uvm_pkg::*;
  import clk_rst_agent_pkg::*;

  //******************************************************************************
  // Includes
  //******************************************************************************
  `include "clk_rst_base_seq.sv"
  `include "clk_rst_mid_sim_rst_seq.sv"

endpackage : clk_rst_seq_pkg