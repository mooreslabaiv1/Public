package rr_agent_pkg;

  //******************************************************************************
  // Imports
  //******************************************************************************
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  //******************************************************************************
  // Includes
  //******************************************************************************
  `include "rr_trans_item.sv"
  `include "rr_monitor.sv"
  `include "rr_driver.sv"
  `include "rr_seqr.sv"
  `include "rr_agent_cov.sv"
  `include "rr_agent_cfg.sv"
  `include "rr_agent.sv"

endpackage : rr_agent_pkg