package requestor_agent_pkg;

  //******************************************************************************
  // Imports
  //******************************************************************************
  import uvm_pkg::*;

  //******************************************************************************
  // Includes
  //******************************************************************************
  `include "requestor_trans_item.sv"
  `include "requestor_monitor.sv"
  `include "requestor_driver.sv"
  `include "requestor_seqr.sv"
  `include "requestor_agent_cov.sv"
  `include "requestor_agent_cfg.sv"
  `include "requestor_agent.sv"

endpackage : requestor_agent_pkg