



    `ifndef SERIALDP_ENV_INC_SV
    `define SERIALDP_ENV_INC_SV
    `include "tb_src.incl"    
    `include "serialDP_env_cfg.sv"
    `include "serialDP_ref_model.sv"
    `include "serialDP_sbd.sv"
    
    `include "serialDP_serial_if_monitor_env_cov.sv"
    `include "serialDP_serial_if_monitor_connect_cov.sv"


    
    `endif // SERIALDP_ENV_INC_SV
    