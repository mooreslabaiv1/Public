package rr_seq_pkg;

  //******************************************************************************
  // Imports
  //******************************************************************************
  import uvm_pkg::*;
  import rr_agent_pkg::*;
  `include "uvm_macros.svh"

  //******************************************************************************
  // Includes
  //******************************************************************************
  `include "rr_base_seq.sv"

endpackage : rr_seq_pkg